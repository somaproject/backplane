library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1A0B844B301B125B842B3FFB100B841B3A1B1A1B840B301B123B888B301B10AB";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"301B137B84AB3FFB100B849B320B120B848B301B12AB846B3FFB100B845B3A0B";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"852B3FFB100B851B3A2B1A2B850B301B13AB84EB302B102B84DB390B190B84CB";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"100B859B321B121B858B301B14BB856B302B102B855B392B192B854B301B147B";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"308B108B860B301B162B85EB302B102B85DB394B194B85CB301B156B85AB3FFB";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"101B869B101B866B3FFB100B865B3A3B1A3B864B301B16EB862B3FFB100B861B";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"A00B100B06D0889B101B1A3A1A2987DB101B879B101B875B101B871B101B86DB";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"374B177B882B36EB165B102D191C809B100B808B101B0B8049E0A00B101B4750";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"882B362B169B880C881B887D20BB300B101B885B36BB12EB884B36FB172B883B";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"3FFB1F0B0B80880C881B887D20BB308B101B885B100B884B100B883B374B100B";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"374B100B884B362B169B883B370B12EB882B364B173B102D191C809B10FB808B";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"1FF7880B190B887B102B0BA0103780B00B80880C881B887D20BB300B101B885B";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"102E103D88348825100C0CA01FF7880B192B20BB101B887B102B100510040C00";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"880B193B885B108B884B100B20BB101B887B102B90C580B4108BCE20B05DA04E";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"101B887B102B0EC010470EA01057A0B8101B4EB0A08B100B0E3010670E101FF7";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"10105020A00B101B4FF0A00B100B0F805040A00B100B0F401077880B194B20BB";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"4BB0A07B100B4F50A07B107B10901087880B131B887B104B1030102010101007";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"108B4ED0A07B106B4E40A07B105B4CB0A07B104B4C10A07B103B46E0A07B101B";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"883B002B882B000B881C001C1290808B0B3B809B0A2B124080BB12204F90A07B";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0C4B80AB0B3B80AB0A2B80DB139010170B311360880D120D887D091D884B032B";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"40BC882B840B881B0A2B14A010470C420B3314608809887B091B80AB0D5B80AB";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"106880C080AB0E6B80AB0D5B80AB0C4B80AB0B3B1550880D121D887D091D883C";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"091B80CB16D0880B109B885B0E6B884B883B882B881B100B887B091B16101057";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"00000000000000000000000000000000000000000000000000001720880A887B";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"AEABB94927ABBBBBBBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"924949B839989266EEE0E0900F9B83A9BB9B7F23AEBAEABBA7F23BBAEBF23AEB";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000001F37B3FEC6BCCCC7B3FB181F3333361ECFFFF731D4924924924926EE56";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
