library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;

library WORK;
use WORK.somabackplane.all;
use work.somabackplane;


library UNISIM;
use UNISIM.VComponents.all;


entity pingdump is
  port (
    CLK      : in  std_logic;
    DOUT      : out std_logic_vector(15 downto 0);
    NEWFRAME : out std_logic);          -- (others => '0')
end pingdump;

architecture Behavioral of pingdump is


  signal netdo   : std_logic_vector(15 downto 0) := (others => '0');
  signal netdop  : std_logic_vector(1 downto 0)  := (others => '0');
  signal netaddr : std_logic_vector(9 downto 0)  := (others => '0');


begin  -- Behavioral

  -- output
  process(CLK)
  begin
    if rising_edge(CLK) then
      DOUT        <= netdo;
      NEWFRAME <= netdop(0);
      netaddr     <= netaddr + 1;
    end if;
  end process;

  RAMB16_S18_inst : RAMB16_S18
    generic map (
      -- Address 0 to 255

      INIT_00  => X"0100A8C054B9014000400200540000450008000100010001FFFFFFFFFFFF0064",
      INIT_01  => X"1312111000000000000EEB6700000000449C24D903000E4BC70200080100A8C0",
      INIT_02  => X"333231302F2E2D2C2B2A292827262524232221201F1E1D1C1B1A191817161514",
      INIT_03  => X"0000000000000000000000000000000000000000000000000000000000003534",
      INIT_04  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F  => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 511
      INIT_10  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F  => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 767
      INIT_20  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F  => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 768 to 1023
      INIT_30  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E  => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F  => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Address 0 to 255
      INITP_00 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Address 768 to 1023
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
      DO       => NETDO,                -- 16-bit Data Output
      DOP      => NETDOP,               -- 2-bit parity Output
      ADDR     => NETADDR,              -- 10-bit Address Input
      CLK      => CLK,                  -- Clock
      DI       => X"0000",
      DIP      => "00",                 -- 2-bit parity Input
      EN       => '1',                  -- RAM Enable Input
      SSR      => '0',                  -- Synchronous Set/Reset Input
      WE       => '0'                   -- Write Enable Input
      );


end Behavioral;
