library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;

library soma;
use soma.somabackplane.all;
use soma.somabackplane;
use soma.all;
library jtag;
use jtag.all;


library network;
use network.all;
library syscon;
use syscon.all;

library UNISIM;
use UNISIM.VComponents.all;

-- for instruction ram for syscontrol

--
entity backplane is
  port (
    CLKIN         : in    std_logic;
    DSPCFG : out std_logic_vector(15 downto 0);
    -- SPI interface
    SPIMOSI       : in    std_logic;
    SPIMISO       : out   std_logic;
    SPICS         : in    std_logic;
    SPICLK        : in    std_logic;
    -- LEDS
    LEDPOWER      : out   std_logic;
    LEDEVENT      : out   std_logic;
    -- NIC interface
    NICFCLK       : out   std_logic;
    NICFDIN       : out   std_logic;
    NICFPROG      : out   std_logic;
    NICSCLK       : out   std_logic;
    NICSIN        : in    std_logic;
    NICSOUT       : out   std_logic;
    NICSCS        : out   std_logic;
    NICDOUT       : out   std_logic_vector(15 downto 0);
    NICNEWFRAME   : out   std_logic;
    NICDIN        : in    std_logic_vector(15 downto 0);
    NICNEXTFRAME  : out   std_logic;
    NICDINEN      : in    std_logic;
    NICIOCLK      : out   std_logic;
    RAMCLKOUT_P   : out   std_logic;
    RAMCLKOUT_N   : out   std_logic;
    RAMCKE        : out   std_logic := '0';
    RAMCAS        : out   std_logic;
    RAMRAS        : out   std_logic;
    RAMCS         : out   std_logic;
    RAMWE         : out   std_logic;
    RAMADDR       : out   std_logic_vector(12 downto 0);
    RAMBA         : out   std_logic_vector(1 downto 0);
    RAMDQSH       : inout std_logic;
    RAMDQSL       : inout std_logic;
    RAMDQ         : inout std_logic_vector(15 downto 0);
    FIBERDEBUGOUT : out   std_logic;
    FIBERDEBUGIN  : in    std_logic;

    -- DeviceLink Serial interfaces
    TXIO_P     : out std_logic_vector(18 downto 0);
    TXIO_N     : out std_logic_vector(18 downto 0);
    RXIO_P     : in  std_logic_vector(18 downto 0);
    RXIO_N     : in  std_logic_vector(18 downto 0)
    );
end backplane;


architecture Behavioral of backplane is

  signal ECYCLE : std_logic := '0';

  signal EARX    : somabackplane.addrarray      := (others => (others => '0'));
  signal EDRX    : somabackplane.dataarray      := (others => (others => '0'));
  signal EDSELRX : std_logic_vector(3 downto 0) := (others => '0');
  signal EATX    : somabackplane.addrarray      := (others => (others => '0'));
  signal EDTX    : std_logic_vector(7 downto 0) := (others => '0');
  signal RESET   : std_logic                    := '0';

  signal lserialboot : std_logic_vector(19 downto 0) := (others => '1');

  signal douta   : std_logic_vector(7 downto 0) := (others => '0');
  signal doutena : std_logic                    := '0';

  signal doutb   : std_logic_vector(7 downto 0) := (others => '0');
  signal doutenb : std_logic                    := '0';


  signal clk, clkint             : std_logic := '0';
  signal clk2x, clk2xint         : std_logic := '0';
  signal clk180, clk180int       : std_logic := '0';
  signal memclkb, memclkbint     : std_logic := '0';
  signal memclk, memclkint       : std_logic := '0';
  signal memclk90, memclk90int   : std_logic := '0';
  signal memclk180, memclk180int : std_logic := '0';
  signal memclk270, memclk270int : std_logic := '0';


  signal nicclkint : std_logic := '0';


-- nic config signals
  signal myip, mybcast : std_logic_vector(31 downto 0) := (others => '0');
  signal mymac         : std_logic_vector(47 downto 0) := (others => '0');

  -- error signals and counters
  signal rxiocrcerr   : std_logic                     := '0';
  signal UNKNOWNETHER : std_logic                     := '0';
  signal UNKNOWNIP    : std_logic                     := '0';
  signal UNKNOWNUDP   : std_logic                     := '0';
  signal UNKNOWNARP   : std_logic                     := '0';
  signal txpktlenen   : std_logic                     := '0';
  signal txpktlen     : std_logic_vector(15 downto 0) := (others => '0');
  signal txchan       : std_logic_vector(2 downto 0)  := (others => '0');
  signal evtrxsuc     : std_logic                     := '0';
  signal evtfifofull  : std_logic                     := '0';


  signal nicnextframeint : std_logic := '0';

  signal locked, locked2 : std_logic                    := '0';
  signal resetint        : std_logic_vector(7 downto 0) := (others => '1');

  signal niciointclk : std_logic                     := '0';
  signal nicdinl     : std_logic_vector(15 downto 0) := (others => '0');
  signal nicdinenl   : std_logic                     := '0';


  signal fiberdebugdest : std_logic_vector(somabackplane.N-1 downto 0) := (others => '0');

  signal fibertxclk, fibertxclkint           : std_logic := '0';
  signal fibertxclkdummy, fibertxclkintdummy : std_logic := '0';

  signal lnicdout     : std_logic_vector(15 downto 0) := (others => '0');
  signal lnicnewframe : std_logic                     := '0';

  signal fiberdebugdebug : std_logic_vector(15 downto 0) := (others => '0');

  signal jtagesenddebug : std_logic_vector(7 downto 0) := (others => '0');

  -- devicelink clocks
  signal clkbittxint, clkbittx       : std_logic := '0';
  signal clkbittx180int, clkbittx180 : std_logic := '0';

  signal clkbitrxint, clkbitrx : std_logic := '0';
  signal clkwordtx       : std_logic := '0';

  signal validint : std_logic_vector(18 downto 0) := (others => '0');

  signal maindcmlocked : std_logic := '0';
  
begin  -- Behavioral


  ---------------------------------------------------------------------------
  -- CLOCKING
  ---------------------------------------------------------------------------

  DCM_BASE_inst : DCM_BASE
    generic map (
      CLKDV_DIVIDE => 2.0,

      CLKFX_DIVIDE          => 1,
      CLKFX_MULTIPLY        => 3,
      CLKIN_DIVIDE_BY_2     => false,
      CLKIN_PERIOD          => 20.0,
      CLKOUT_PHASE_SHIFT    => "NONE",
      CLK_FEEDBACK          => "1X",
      DCM_AUTOCALIBRATION   => true,
      DFS_FREQUENCY_MODE    => "LOW",
      DLL_FREQUENCY_MODE    => "LOW",
      DUTY_CYCLE_CORRECTION => true,
      STARTUP_WAIT          => true)
    port map (
      CLK0                  => clkint,      -- 0 degree DCM CLK ouptput
      CLK2x                 => clk2xint,
      CLKFX                 => memclkbint,  -- DCM CLK synthesis out (M/D)
      CLKFB                 => clk,
      CLK180                => clk180int,
      CLK90                 => niciointclk,
      CLKIN                 => CLKIN,
      LOCKED                => locked,
      RST                   => '0'          -- DCM asynchronous reset input
      );

  clk_bufg : BUFG
    port map (
      O => clk,
      I => clkint);

  clk180_bufg : BUFG
    port map (
      I => clk180int,
      O => clk180);

  clk2x_bufg : BUFG
    port map (
      I => clk2xint,
      O => clk2x);

  memclkb_bufg : BUFG
    port map (
      O => memclkb,
      I => memclkbint);

  process(CLK)
  begin
    if rising_edge(CLK) then
      resetint <= resetint(6 downto 0) & (not locked);
    end if;
  end process;


  DCM_BASE_inst2 : DCM_BASE
    generic map (
      CLKDV_DIVIDE => 2.0,

      CLKIN_DIVIDE_BY_2     => false,
      CLKIN_PERIOD          => 6.0,
      CLKOUT_PHASE_SHIFT    => "NONE",
      CLK_FEEDBACK          => "1X",
      DCM_AUTOCALIBRATION   => true,
      DCM_PERFORMANCE_MODE  => "MAX_SPEED",
      DESKEW_ADJUST         => "SYSTEM_SYNCHRONOUS",
      DFS_FREQUENCY_MODE    => "LOW",
      DLL_FREQUENCY_MODE    => "LOW",
      DUTY_CYCLE_CORRECTION => true,
      STARTUP_WAIT          => false)
    port map (
      CLK0                  => memclkint,
      CLK180                => memclk180int,
      CLK270                => memclk270int,
      CLK90                 => memclk90int,
      CLKFB                 => memclk,
      CLKIN                 => memclkb,
      LOCKED                => locked2,
      RST                   => resetint(7)

      );

  RESET <= not locked2;

  memclk_bufg : BUFG
    port map (
      O => memclk,
      I => memclkint);

  memclk90_bufg : BUFG
    port map (
      O => memclk90,
      I => memclk90int);

  memclk180_bufg : BUFG
    port map (
      O => memclk180,
      I => memclk180int);

  memclk270_bufg : BUFG
    port map (
      O => memclk270,
      I => memclk270int);

  TXIO_obufds : OBUFDS
    generic map (
      IOSTANDARD => "DEFAULT")
    port map (
      O          => RAMCLKOUT_P,
      OB         => RAMCLKOUT_N,
      I          => memclk270
      );

  eventrouter_inst : entity soma.eventrouter
    port map (
      CLK     => clk,
      ECYCLE  => ECYCLE,
      EARX    => EARX,
      EDRX    => EDRX,
      EDSELRX => EDSELRX,
      EATX    => EATX,
      EDTX    => EDTX);

  timer_inst      : entity soma.timer
    port map (
      CLK         => clk,
      ECYCLe      => ECYCLE,
      EARX        => EARX(0),
      EDRX        => EDRX(0),
      EDSELRX     => EDSELRX,
      EATX        => EATX(0),
      EDTX        => EDTX);
  -- init syscontrol with the ram values so that we can properly sim
  syscontrol_inst : entity syscon.syscontrol
    generic map (
      RAM_INIT_00 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_00,
      RAM_INIT_01 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_01,
      RAM_INIT_02 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_02,
      RAM_INIT_03 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_03,
      RAM_INIT_04 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_04,
      RAM_INIT_05 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_05,
      RAM_INIT_06 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_06,
      RAM_INIT_07 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_07,
      RAM_INIT_08 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_08,
      RAM_INIT_09 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_09,
      RAM_INIT_0A => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0A,
      RAM_INIT_0B => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0B,
      RAM_INIT_0C => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0C,
      RAM_INIT_0D => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0D,
      RAM_INIT_0E => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0E,
      RAM_INIT_0F => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_0F,

      RAM_INIT_10 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_10,
      RAM_INIT_11 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_11,
      RAM_INIT_12 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_12,
      RAM_INIT_13 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_13,
      RAM_INIT_14 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_14,
      RAM_INIT_15 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_15,
      RAM_INIT_16 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_16,
      RAM_INIT_17 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_17,
      RAM_INIT_18 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_18,
      RAM_INIT_19 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_19,
      RAM_INIT_1A => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1A,
      RAM_INIT_1B => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1B,
      RAM_INIT_1C => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1C,
      RAM_INIT_1D => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1D,
      RAM_INIT_1E => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1E,
      RAM_INIT_1F => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_1F,

      RAM_INIT_20 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_20,
      RAM_INIT_21 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_21,
      RAM_INIT_22 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_22,
      RAM_INIT_23 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_23,
      RAM_INIT_24 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_24,
      RAM_INIT_25 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_25,
      RAM_INIT_26 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_26,
      RAM_INIT_27 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_27,
      RAM_INIT_28 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_28,
      RAM_INIT_29 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_29,
      RAM_INIT_2A => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2A,
      RAM_INIT_2B => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2B,
      RAM_INIT_2C => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2C,
      RAM_INIT_2D => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2D,
      RAM_INIT_2E => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2E,
      RAM_INIT_2F => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_2F,

      RAM_INIT_30 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_30,
      RAM_INIT_31 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_31,
      RAM_INIT_32 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_32,
      RAM_INIT_33 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_33,
      RAM_INIT_34 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_34,
      RAM_INIT_35 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_35,
      RAM_INIT_36 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_36,
      RAM_INIT_37 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_37,
      RAM_INIT_38 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_38,
      RAM_INIT_39 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_39,
      RAM_INIT_3A => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3A,
      RAM_INIT_3B => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3B,
      RAM_INIT_3C => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3C,
      RAM_INIT_3D => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3D,
      RAM_INIT_3E => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3E,
      RAM_INIT_3F => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INIT_3F,

      RAM_INITP_00 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_00,
      RAM_INITP_01 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_01,
      RAM_INITP_02 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_02,
      RAM_INITP_03 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_03,
      RAM_INITP_04 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_04,
      RAM_INITP_05 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_05,
      RAM_INITP_06 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_06,
      RAM_INITP_07 => work.backplane_mem_pkg.syscontrol_inst_instruction_ram_INITP_07)
    port map (
      CLK          => clk,
      CLK2X        => clk2x,
      RESET        => RESET,
      ECYCLe       => ECYCLE,
      EARX         => EARX(1),
      EDRX         => EDRX(1),
      EDSELRX      => EDSELRX,
      EATX         => EATX(1),
      EDTX         => EDTX,
      SEROUT       => lserialboot);

  bootstore_inst : entity soma.bootstore
    generic map (
      DEVICE  => X"02")
    port map (
      CLK     => clk,
      CLKHI   => memclk,
      RESET   => RESET,
      ECYCLE  => ECYCLE,
      EARX    => EARX(2),
      EDRX    => EDRX(2),
      EDSELRX => EDSELRX,
      EATX    => EATX(2),
      EDTX    => EDTX,
      SPIMOSI => SPIMOSI,
      SPIMISO => SPIMISO,
      SPICS   => SPICS,
      SPICLK  => SPICLK);

  bootdeserialize_inst : entity soma.bootdeserialize
    port map (
      CLK   => clk,
      SERIN => lserialboot(0),
      FPROG => NICFPROG,
      FCLK  => NICFCLK,
      FDIN  => NICFDIN);

  DSPCFG <= lserialboot(19 downto 4);


  LEDPOWER <= lserialboot(0);
  LEDEVENT <= jtagesenddebug(1);

  jtagsend_inst : entity jtag.jtagesend
    generic map (
      JTAG_CHAIN => 1)
    port map (
      CLK        => clk,
      ECYCLE     => ecycle,
      EARX       => earx(7),
      EDRX       => edrx(7),
      EDSELRX    => edselrx,
      DEBUG      => jtagesenddebug);

  jtagreceive_inst : entity jtag.jtagereceive
    generic map (
      JTAG_CHAIN_MASK => 2,
      JTAG_CHAIN_OUT  => 3 )
    port map (
      CLK             => clk,
      ECYCLE          => ecycle,
      EDTX            => edtx,
      EATX            => eatx(7),
      DEBUG           => open);

  DCM_fibertx_inst : DCM_BASE
    generic map (
      CLKFX_DIVIDE   => 5,
      CLKFX_MULTIPLY => 8,
      STARTUP_WAIT   => true)
    port map (
      CLKFX          => fibertxclkint,
      CLKIN          => clk,
      CLK0           => fibertxclkintdummy,
      CLKFB          => fibertxclkdummy,
      LOCKED         => open,
      RST            => '0'             -- DCM asynchronous reset input
      );

  clk_fibertx_bufg : BUFG
    port map (
      O => fibertxclk,
      I => fibertxclkint);

  clk_fibertxdummy_bufg : BUFG
    port map (
      O => fibertxclkdummy,
      I => fibertxclkintdummy);

  fiberdebug_inst : entity soma.fiberdebug
    generic map (
      DEVICE    => X"4C")
    port map (
      CLK       => CLK,
      TXCLK     => fibertxclk,
      RESET     => reset,
      ECYCLE    => ecycle,
      EARXA     => earx(70),
      EDRXA     => edrx(70),
      EDSELRXA  => edselrx,
      EARXB     => earx(71),
      EDRXB     => edrx(71),
      EDSELRXB  => edselrx,
      EATX      => eatx(70),
      EDTX      => edtx,
      EADDRDEST => fiberdebugdest,
      FIBERIN   => FIBERDEBUGIN,
      FIBEROUT  => FIBERDEBUGOUT,
      DEBUG     => fiberdebugdebug);


  fakedata1 : entity work.fakedata
    port map (
      clk    => clk,
      DOUT   => douta,
      DOUTEN => doutena,
      ECYCLE => ecycle);

  -- dummy
  process(clk)
    variable blinkcnt : std_logic_vector(21 downto 0)
               := (others => '0');
  begin
    if rising_edge(clk) then
      blinkcnt := blinkcnt + 1;

    end if;
  end process;

-- NETCLK <= clk;



-- myip <= X"0A000002";                 -- 10.0.0.2
--   mybcast <= X"FFFFFFFF";            -- 10.255.255.255

-- mymac <= X"00ADBEEF1234";

  fiberdebugdest(3) <= '1';
  network_inst : entity network.network
    port map (
      CLK       => CLK,
      MEMCLK    => memclk,
      MEMCLK90  => memclk90,
      MEMCLK180 => memclk180,
      MEMCLK270 => memclk270,
      RESET     => RESET,
      -- config
      MYIP      => MYIP,
      MYMAC     => mymac,
      MYBCAST   => mybcast,

      -- input
      NICNEXTFRAME => NICNEXTFRAME,
      NICDINEN     => nicdinenl,
      NICDIN       => nicdinl,
      -- output
      NICDOUT      => lNICDOUT,
      NICNEWFRAME  => lNICNEWFRAME,
      NICIOCLK     => open,             --NICIOCLK,
      -- event bus
      ECYCLE       => ecycle,
      EARX         => earx(3),
      EDRX         => edrx(3),
      EDSELRX      => edselrx,
      EATX         => eatx(3),
      EDTX         => edtx,

      -- data bus
      DIENA => doutena,
      DIENB => '0',
      DINA  => douta,
      DINB  => X"00",

      -- memory interface
      RAMCKE  => RAMCKE,
      RAMCAS  => RAMCAS,
      RAMRAS  => RAMRAS,
      RAMCS   => RAMCS,
      RAMWE   => RAMWE,
      RAMADDR => RAMADDR,
      RAMBA   => RAMBA,
      RAMDQSH => RAMDQSH,
      RAMDQSL => RAMDQSL,
      RAMDQ   => RAMDQ,

      -- counters
      RXIOCRCERR   => rxiocrcerr,
      UNKNOWNETHER => unknownether,
      UNKNOWNIP    => unknownip,
      UNKNOWNUDP   => unknownudp,
      UNKNOWNARP   => unknownarp,
      TXPKTLENEN   => txpktlenen,
      TXPKTLEN     => txpktlen,
      TXCHAN       => txchan,
      EVTRXSUC     => evtrxsuc,
      EVTFIFOFULL  => evtfifofull

      );

  netcontrol_inst : entity soma.netcontrol
    generic map (
      DEVICE      => X"04"
--       RAM_INIT_00 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_00,
--       RAM_INIT_01 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_01,
--       RAM_INIT_02 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_02,
--       RAM_INIT_03 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_03,
--       RAM_INIT_04 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_04,
--       RAM_INIT_05 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_05,
--       RAM_INIT_06 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_06,
--       RAM_INIT_07 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_07,
--       RAM_INIT_08 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_08,
--       RAM_INIT_09 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_09,
--       RAM_INIT_0A => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0A,
--       RAM_INIT_0B => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0B,
--       RAM_INIT_0C => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0C,
--       RAM_INIT_0D => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0D,
--       RAM_INIT_0E => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0E,
--       RAM_INIT_0F => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_0F,

--       RAM_INIT_10 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_10,
--       RAM_INIT_11 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_11,
--       RAM_INIT_12 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_12,
--       RAM_INIT_13 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_13,
--       RAM_INIT_14 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_14,
--       RAM_INIT_15 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_15,
--       RAM_INIT_16 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_16,
--       RAM_INIT_17 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_17,
--       RAM_INIT_18 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_18,
--       RAM_INIT_19 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_19,
--       RAM_INIT_1A => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1A,
--       RAM_INIT_1B => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1B,
--       RAM_INIT_1C => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1C,
--       RAM_INIT_1D => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1D,
--       RAM_INIT_1E => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1E,
--       RAM_INIT_1F => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_1F,

--       RAM_INIT_20 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_20,
--       RAM_INIT_21 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_21,
--       RAM_INIT_22 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_22,
--       RAM_INIT_23 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_23,
--       RAM_INIT_24 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_24,
--       RAM_INIT_25 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_25,
--       RAM_INIT_26 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_26,
--       RAM_INIT_27 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_27,
--       RAM_INIT_28 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_28,
--       RAM_INIT_29 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_29,
--       RAM_INIT_2A => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2A,
--       RAM_INIT_2B => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2B,
--       RAM_INIT_2C => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2C,
--       RAM_INIT_2D => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2D,
--       RAM_INIT_2E => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2E,
--       RAM_INIT_2F => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_2F,

--       RAM_INIT_30 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_30,
--       RAM_INIT_31 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_31,
--       RAM_INIT_32 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_32,
--       RAM_INIT_33 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_33,
--       RAM_INIT_34 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_34,
--       RAM_INIT_35 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_35,
--       RAM_INIT_36 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_36,
--       RAM_INIT_37 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_37,
--       RAM_INIT_38 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_38,
--       RAM_INIT_39 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_39,
--       RAM_INIT_3A => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3A,
--       RAM_INIT_3B => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3B,
--       RAM_INIT_3C => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3C,
--       RAM_INIT_3D => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3D,
--       RAM_INIT_3E => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3E,
--       RAM_INIT_3F => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INIT_3F,

--       RAM_INITP_00 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_00,
--       RAM_INITP_01 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_01,
--       RAM_INITP_02 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_02,
--       RAM_INITP_03 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_03,
--       RAM_INITP_04 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_04,
--       RAM_INITP_05 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_05,
--       RAM_INITP_06 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_06,
--       RAM_INITP_07 => work.backplane_mem_pkg.netcontrol_inst_instruction_ram_INITP_07)
      )
    port map (
      CLK          => CLK,
      CLK2X        => CLK2X,
      RESET        => RESET,
      -- standard event-bus interface
      ECYCLE       => ECYCLE,
      EDTX         => EDTX,
      EATX         => EATX(4),
      EARX         => EARX(4),
      EDRX         => EDRX(4),
      EDSELRX      => EDSELRX,
      -- tx counter input
      TXPKTLENEN   => txpktlenen,
      TXPKTLEN     => txpktlen,
      TXCHAN       => txchan,
      -- other counters
      RXIOCRCERR   => rxiocrcerr,
      UNKNOWNETHER => unknownether,
      UNKNOWNIP    => unknownip,
      UNKNOWNARP   => unknownarp,
      UNKNOWNUDP   => unknownudp,
      EVTRXSUC     => evtrxsuc,
      EVTFIFOFULL  => evtfifofull,
      -- output network control settings
      MYMAC        => mymac,
      MYBCAST      => mybcast,
      MYIP         => myip,
      -- NIC interface
      NICSOUT      => NICSOUT,
      NICSIN       => NICSIN,
      NICSCLK      => NICSCLK,
      NICSCS       => NICSCS
      );


  NICIOCLK <= clk;

  process(niciointclk)
  begin

    if rising_edge(niciointclk) then
      nicdinenl <= NICDINEN;
      nicdinl   <= NICDIN;

    end if;

  end process;

  process(CLK)
  begin
    if rising_edge(CLK) then
      NICDOUT     <= lnicdout;
      NICNEWFRAME <= lnicnewframe;

    end if;
  end process;


    devicelinkclk_inst : entity work.devicelinkclk
    port map (
      CLKIN       => CLKIN,
      CLKBITTX    => clkbittx,
      CLKBITTX180 => clkbittx180,
      CLKBITRX    => clkbitrx,
      CLKWORDTX   => clkwordtx,
      STARTUPDONE => maindcmlocked);
  
  -- instantiate devices

   devicelinks : for i in 0 to 15 generate
     dl        : entity work.linktester
       port map (
         CLK       => clk,
         RXBITCLK  => clkbitrx,
         TXHBITCLK => clkbittx,
         TXWORDCLK => clkwordtx,
         RESET     => RESET,
         TXIO_P    => TXIO_P(i),
         TXIO_N    => TXIO_N(i),
         RXIO_P    => RXIO_P(i),
         RXIO_N    => RXIO_N(i),
         VALID     => validint(i));

   end generate devicelinks;


end Behavioral;
