library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;

library WORK;
use WORK.somabackplane.all;
use work.somabackplane;



entity syscontroltest is
  
end syscontroltest;


architecture Behavioral of syscontroltest is

begin  -- Behavioral

  

end Behavioral;
