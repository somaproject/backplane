
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package somabackplane is

  type dataarray is array(39 downto 0) of std_logic_vector(7 downto 0); 
  
end somabackplane;


package body somabackplane is

 
end somabackplane;
