library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1929844930091FA9842930291029841939091909840930091F79888930091DE9";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"301910B984A93FF91009849932091209848930091FE984693029102984593929";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"101985D9101985991019855910198519101984E93029102984D93949194984C9";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"101987D9101987991019875910198719101986D9101986991019865910198619";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"1659102B191A809910098089101908C04720A00910194490A009100904108899";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"8819887B209930091019885936B912E9884936F91729883937491779882936E9";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"8819887B2099308910198859100988491009883937491009882936291699880A";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"16998839370912E9882936491739102B191A809910F980893FF91F0908C0880A";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"102908E0103780B008C0880A8819887B20993009101988593749100988493629";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"100A09E01FF78809192920991019887910291005100409401FF7880919098879";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"88491009209910198879102990A580941089CB60B05BA04C102C103B88348825";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"10470BE01057A09810194BF0A08910090B7010670B501FF78809193988591089";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"4D30A00910090CC04D80A00910090C8010778809194920991019887910290C00";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"A07910790DD0108788091319887910490D700D600D50100710104D60A0091019";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"4B80A079105949F0A07910494950A07910394420A079101948F0A07910094C90";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"881A001A0FD010470C420B330F9010170B310F604CD0A07910894C10A0791069";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"0D5980A90C4980A90B3910A0880B120B887B091B884903298839002988290009";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"00000000000000000000000000000000000011601057106880C080A90E6980A9";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"BAEABBA7F23BBAEBF23AEBAEABB94927BBBBBBBBBBBBBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"F60614924924924926EE56924949B839989266EEE0E0900F9B83A9BB9B7F23AE";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"00000000000000000000000000000000000000000000000000001AF3331ECFFF";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1416844630061C4684263FF61006841633161316840630061C16888630061B96";
		constant netcontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"30061D5684A63FF61006849634061406848630061C8684663FF6100684563416";
		constant netcontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"101685D6101685961016855610168516101684E63FF6100684D63306130684C6";
		constant netcontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"140487D6101687961016875610168716101686D6101686961016865610168616";
		constant netcontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"A01610164660A016100604A08806130688728827883600370046042088951015";
		constant netcontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"48D0A01610464AD0A01610764A20A01610664860A016103647C0A016102646E0";
		constant netcontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"1016000706D010118006804680368026801610064B70A0161FF649A0A0161056";
		constant netcontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"100680268016101607B010210790100147A0A07600373016123607204730A076";
		constant netcontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"10968016101608C0104108A048B0A07610160007085010318006804610168036";
		constant netcontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"09F04A00A0361006A063101609903F0310031051800680468036311614068026";
		constant netcontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"A076101600070AC010718006804612068036100680261086801610160A101061";
		constant netcontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"4430A0651015000644B0A00510150B8010000B601FF18806887610760B104B20";
		constant netcontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"406A40694068820688160A26887709170C70C06682060A260C30100110100C00";
		constant netcontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"0DF08005091280450D5580350C4580250B3580150A250D408804884A88398828";
		constant netcontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"BE664E94B6FFE49249249249249EFFDEBBBBBBBBBBBBBAEBAEBAEBAEBAEBAEBA";
		constant netcontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"0000000000000000733331FFFECC78694B499BE52DBEEEE65226AFEBB994B6FB";
		constant netcontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
end backplane_mem_pkg;
