library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1A0B844B301B12CB842B3FFB100B841B3A1B1A1B840B301B12AB888B301B111B";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"301B13EB84AB3FFB100B849B320B120B848B301B131B846B3FFB100B845B3A0B";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"852B3FFB100B851B322B122B850B301B141B84EB302B102B84DB390B190B84CB";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"100B859B321B121B858B301B150B856B302B102B855B392B192B854B301B14CB";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"308B108B860B301B167B85EB302B102B85DB394B194B85CB301B15BB85AB3FFB";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"868B301B178B866B3FFB100B865B3A3B1A3B864B301B173B862B3FFB100B861B";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"87DB101B879B101B875B101B871B101B86DB101B86AB3FFB100B869B3A2B1A2B";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"809B100B808B101B0BF04A50A00B101B47C0A00B100B0740889B101B1A3A1A29";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"300B101B885B36BB12EB884B36FB172B883B374B177B882B36EB165B102D191C";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"308B101B885B100B884B100B883B374B100B882B362B169B880C881B887D20BB";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"12EB882B364B173B102D191C809B10FB808B3FFB1F0B0BF0880C881B887D20BB";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"80B00BF0880C881B887D20BB300B101B885B374B100B884B362B169B883B370B";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"880B192B20BB101B887B102B100510040C701FF7880B190B887B102B0C101037";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"101B887B102B90C580B4108BCE90B05DA04E102E103D88348825100C0D101FF7";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"A0B8101B4F20A08B100B0EA010670E801FF7880B193B885B108B884B100B20BB";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"0FF050B0A00B100B0FB01077880B194B20BB101B887B102B0F3010470F101057";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"1087880B131B887B104B10A010901080100710105090A00B101B5060A00B100B";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"4D20A07B104B4C80A07B103B4750A07B101B4C20A07B100B4FC0A07B107B1100";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"808B0B3B809B0A2B12B080BB12905000A07B108B4F40A07B106B4EB0A07B105B";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"10170B3113D0880D120D887D091D884B032B883B002B882B000B881C001C1300";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"14F010470C420B3314B0880B122B882B051B051B881B050B050B887B091B1400";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0D5B80AB0C4B80AB0B3B15A0880D121D887D091D883C40BC882B840B881B0A2B";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"885B0E6B884B883B882B881B100B887B091B16601057106880C080AB0E6B80AB";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0D5B80AB0C4B80AB0B3B80AB0A2B80DB1770880A887B091B80CB1720880B109B";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000018408809887B091B80AB";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"EE5249EAEEEEEEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"526E0E662499BBB8382403E6E0EA6EE6DFC8EBAEBAAEE9FC8EEEBAFC8EBAEBAA";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"33337CDECFFB1AF3331ECFEC607BFFF187B3FFFDCC75249249249249BB95A492";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"00000000000000000000000000000000000000000000000000000000000001F3";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
