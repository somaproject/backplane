library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

entity bitcnt is
  port (
    CLK   : in  std_logic;
    DIN   : in  std_logic_vector(95 downto 0);
    DOUT  : out std_logic_vector(6 downto 0);
    START : in  std_logic;
    DONE  : out std_logic
    );
end bitcnt;

architecture Behavioral of bitcnt is
  signal do : std_logic_vector(31 downto 0) := (others => '0');
  signal s1 : std_logic_vector(19 downto 0) := (others => '0');
  signal s2 : std_logic_vector(11 downto 0) := (others => '0');

  signal w1, w2, w3 : std_logic := '0';


begin  -- Behavioral

  darray : for i in 0 to 3 generate
    mem  : RAMB16_S4_S4
      generic map (
        SIM_COLLISION_CHECK => "NONE",
        INIT_00             => X"6554544354434332544343324332322154434332433232214332322132212110",
        INIT_01             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_02             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_03             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_04             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_05             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_06             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_07             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_08             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_09             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_0A             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_0B             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_0C             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_0D             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_0E             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_0F             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_10             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_11             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_12             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_13             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_14             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_15             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_16             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_17             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_18             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_19             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_1A             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_1B             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_1C             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_1D             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_1E             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_1F             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_20             => X"7665655465545443655454435443433265545443544343325443433243323221",
        INIT_21             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_22             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_23             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_24             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_25             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_26             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_27             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_28             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_29             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_2A             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_2B             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_2C             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_2D             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_2E             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_2F             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_30             => X"8776766576656554766565546554544376656554655454436554544354434332",
        INIT_31             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_32             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_33             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_34             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_35             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_36             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_37             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_38             => X"9887877687767665877676657665655487767665766565547665655465545443",
        INIT_39             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_3A             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_3B             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_3C             => X"A998988798878776988787768776766598878776877676658776766576656554",
        INIT_3D             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_3E             => X"BAA9A998A9989887A998988798878776A9989887988787769887877687767665",
        INIT_3F             => X"CBBABAA9BAA9A998BAA9A998A9989887BAA9A998A9989887A998988798878776"
        )
      port map (
        WEA   => '0',
        ENA   => '1',
        SSRA  => '0',
        CLKA  => CLK,
        ADDRA => DIN(24*i+11 downto 24*i),
        ADDRB => DIN(24*i+23 downto 24*i + 12),
        DIA   => "0000",
        DOA   => do(8*i+3 downto 8*i),
        WEB   => '0',
        ENB   => '1',
        SSRB  => '0',
        CLKB  => CLK,
        DIB   => "0000",
        DOB   => do(8*i+7 downto 8*i+4));

    process (CLK)
    begin
      if rising_edge(CLK) then
        s1(5*i +4 downto 5*i) <= ('0' & do(8*i+3 downto 8*i))
                                 + ('0' & do(8*i+7 downto 8*i+4));
      end if;
    end process;
  end generate darray;

  darray2 : for i in 0 to 1 generate
    process (CLK)
    begin
      if rising_edge(CLK) then
        s2(6*i +5 downto 6*i) <= ('0' & s1(10*i +4 downto 10*i)) +
                                 ('0' & s1(10*i +9 downto 10*i+5));
      end if;
    end process;
  end generate darray2;

  main : process(CLK)
  begin
    if rising_edge(CLK) then
      DOUT <= ('0' & s2(5 downto 0)) + ('0' & s2(11 downto 6));
      w1 <= START;
      w2 <= W1;
      W3 <= W2;
      DONE <= w3; 
    end if;
  end process main;
end Behavioral;
