library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"120B844B301B121B842B3FFB100B841B3A0B1A0B840B301B11CB888B301B103B";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"301B131B84AB302B102B849B390B190B848B301B12EB846B3FFB100B845B320B";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"852B302B102B851B392B192B850B301B13EB84EB3FFB100B84DB3A2B1A2B84CB";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"102B859B394B194B858B301B144B856B3FFB100B855B3A1B1A1B854B301B142B";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"3A3B1A3B860B301B15CB85EB3FFB100B85DB308B108B85CB301B150B85AB302B";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"879B101B875B101B871B101B86DB101B869B101B865B101B862B3FFB100B861B";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"808B101B0B104970A00B101B46E0A00B100B0660889B101B1A3A1A2987DB101B";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"885B36BB12EB884B36FB172B883B374B177B882B36EB165B102D191C809B100B";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"885B100B884B100B883B374B100B882B362B169B880C881B887D20BB300B101B";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"364B173B102D191C809B10FB808B3FFB1F0B0B10880C881B887D20BB308B101B";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"880C881B887D20BB300B101B885B374B100B884B362B169B883B370B12EB882B";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"20BB101B887B102B100510040B901FF7880B190B887B102B0B30103780B00B10";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"102B90C580B4108BCDB0B05DA04E102E103D88348825100C0C301FF7880B192B";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"4E40A08B100B0DC010670DA01FF7880B193B885B108B884B100B20BB101B887B";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"A00B100B0ED01077880B194B20BB101B887B102B0E5010470E301057A0B8101B";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"131B887B104B0FC00FB00FA0100710104FB0A00B101B4F80A00B100B0F104FD0";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"104B4BA0A07B103B4670A07B101B4B40A07B100B4EE0A07B107B10201087880B";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"808B0B3B809B0A2B11B04F20A07B108B4E60A07B106B4DD0A07B105B4C40A07B";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"10170B3112D0880D120D887D091D884B032B883B002B882B000B881C001C1200";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0C420B3313D08809887B091B80AB0D5B80AB0C4B80AB0B3B80AB0A2B80DB1300";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"14F01057106880C080AB0E6B80AB0D5B80AB0C4B80AB0B3B143080BB14101047";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"880A887B091B80CB15B0880B109B885B0E6B884B883B882B881B100B887B091B";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000001600";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"EBAEBAAEE5249EAEEEEEEEEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"B95A492526E0E662499BBB8382403E6E0EA6EE6DFC8EBAEBAAEE9FC8EEEBAFC8";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000000000000001F37B3FEC6BCCCC7607CCCCCD87B3FFFDCC5249249249249B";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1416844630061C4684263FF61006841633161316840630061C16888630061B96";
		constant netcontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"30061D5684A63FF61006849634061406848630061C8684663FF6100684563416";
		constant netcontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"101685D6101685961016855610168516101684E63FF6100684D63306130684C6";
		constant netcontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"140487D6101687961016875610168716101686D6101686961016865610168616";
		constant netcontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"A01610164660A016100604A08806130688728827883600370046042088951015";
		constant netcontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"48D0A01610464AD0A01610764A20A01610664860A016103647C0A016102646E0";
		constant netcontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"1016000706D010118006804680368026801610064B70A0161FF649A0A0161056";
		constant netcontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"100680268016101607B010210790100147A0A07600373016123607204730A076";
		constant netcontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"10968016101608C0104108A048B0A07610160007085010318006804610168036";
		constant netcontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"09F04A00A0361006A063101609903F0310031051800680468036311614068026";
		constant netcontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"A076101600070AC010718006804612068036100680261086801610160A101061";
		constant netcontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"4430A0651015000644B0A00510150B8010000B601FF18806887610760B104B20";
		constant netcontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"406A40694068820688160A26887709170C70C06682060A260C30100110100C00";
		constant netcontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"0DF08005091280450D5580350C4580250B3580150A250D408804884A88398828";
		constant netcontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"BE664E94B6FFE49249249249249EFFDEBBBBBBBBBBBBBAEBAEBAEBAEBAEBAEBA";
		constant netcontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"0000000000000000733331FFFECC78694B499BE52DBEEEE65226AFEBB994B6FB";
		constant netcontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
end backplane_mem_pkg;
