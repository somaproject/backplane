library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"180984493019119984293FF910098419320912098409301910C9888930091F39";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"3019121984A9302910298499390919098489301911E984693FF9100984593809";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"8529302910298519392919298509301912B984E93FF9100984D93829182984C9";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"102985993949194985893019131985693FF910098559381918198549301912F9";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"875910198719101986D9101986991019865910198619101985D9101985A93029";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"808910190A104870A009101945E0A009100905608899101987D9101987991019";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"885936B912E9884936F91729883937491779882936E91659102B191A80991009";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"8859100988491009883937491009882936291699880A8819887B209930091019";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"36491739102B191A809910F980893FF91F090A10880A8819887B209930891019";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"880A8819887B2099300910198859374910098849362916998839370912E98829";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"2099101988791029100510040A901FF788091909887910290A30103780B00A10";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"102990A580941089CCB0B05BA04C102C103B88348825100A0B301FF788091929";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"4D40A08910090CC010670CA01FF7880919398859108988491009209910198879";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"A00910090DD010778809194920991019887910290D5010470D301057A0981019";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"1319887910490EC00EB00EA0100710104EB0A00910194E80A00910090E104ED0";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"10494AA0A07910394570A07910194A40A07910094DE0A07910790F2010878809";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"88290009881A001A10B04E20A07910894D60A07910694CD0A07910594B40A079";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"10170B3111D080890B3980990A291180880B120B887B091B8849032988390029";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"80B912E010470C420B3312A080C080A90D5980A90C4980A90B3980A90A291200";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"00000000000013C01057106880C080A90E6980A90D5980A90C4980A90B391300";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"EEEBAFC8EBAEBAAEE5249EEEEEEEEEEEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"9249249BB95A492526E0E662499BBB8382403E6E0EA6EE6DFC8EBAEBAAEE9FC8";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000000000000000000000000000000001AF3331D81F33318731ECFFFF524924";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1416844630061C4684263FF61006841633161316840630061C16888630061B96";
		constant netcontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"30061D5684A63FF61006849634061406848630061C8684663FF6100684563416";
		constant netcontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"101685D6101685961016855610168516101684E63FF6100684D63306130684C6";
		constant netcontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"140487D6101687961016875610168716101686D6101686961016865610168616";
		constant netcontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"A01610164660A016100604A08806130688728827883600370046042088951015";
		constant netcontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"48D0A01610464AD0A01610764A20A01610664860A016103647C0A016102646E0";
		constant netcontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"1016000706D010118006804680368026801610064B70A0161FF649A0A0161056";
		constant netcontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"100680268016101607B010210790100147A0A07600373016123607204730A076";
		constant netcontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"10968016101608C0104108A048B0A07610160007085010318006804610168036";
		constant netcontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"09F04A00A0361006A063101609903F0310031051800680468036311614068026";
		constant netcontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"A076101600070AC010718006804612068036100680261086801610160A101061";
		constant netcontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"4430A0651015000644B0A00510150B8010000B601FF18806887610760B104B20";
		constant netcontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"406A40694068820688160A26887709170C70C06682060A260C30100110100C00";
		constant netcontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"0DF08005091280450D5580350C4580250B3580150A250D408804884A88398828";
		constant netcontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"BE664E94B6FFE49249249249249EFFDEBBBBBBBBBBBBBAEBAEBAEBAEBAEBAEBA";
		constant netcontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"0000000000000000733331FFFECC78694B499BE52DBEEEE65226AFEBB994B6FB";
		constant netcontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant netcontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
end backplane_mem_pkg;
