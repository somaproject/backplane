library ieee;
use ieee.std_logic_1164;
package backplane_mem_pkg is
		constant syscontrol_inst_instruction_ram_INIT_00 : bit_vector(0 to 255) := X"1A0C844C301C12CC842C3FFC100C841C3A1C1A1C840C301C12AC888C301C111C";
		constant syscontrol_inst_instruction_ram_INIT_01 : bit_vector(0 to 255) := X"301C13EC84AC3FFC100C849C320C120C848C301C131C846C3FFC100C845C3A0C";
		constant syscontrol_inst_instruction_ram_INIT_02 : bit_vector(0 to 255) := X"852C3FFC100C851C322C122C850C301C141C84EC302C102C84DC390C190C84CC";
		constant syscontrol_inst_instruction_ram_INIT_03 : bit_vector(0 to 255) := X"100C859C321C121C858C301C152C856C302C102C855C392C192C854C301C14EC";
		constant syscontrol_inst_instruction_ram_INIT_04 : bit_vector(0 to 255) := X"308C108C860C301C16BC85EC302C102C85DC394C194C85CC301C15FC85AC3FFC";
		constant syscontrol_inst_instruction_ram_INIT_05 : bit_vector(0 to 255) := X"868C301C17CC866C3FFC100C865C3A3C1A3C864C301C177C862C3FFC100C861C";
		constant syscontrol_inst_instruction_ram_INIT_06 : bit_vector(0 to 255) := X"87DC101C879C101C875C101C871C101C86DC101C86AC3FFC100C869C3A2C1A2C";
		constant syscontrol_inst_instruction_ram_INIT_07 : bit_vector(0 to 255) := X"809C100C808C101C0BF04A50A00C101C47C0A00C100C0740889C101C1A3A1A29";
		constant syscontrol_inst_instruction_ram_INIT_08 : bit_vector(0 to 255) := X"300C101C885C36BC12EC884C36FC172C883C374C177C882C36EC165C102E191D";
		constant syscontrol_inst_instruction_ram_INIT_09 : bit_vector(0 to 255) := X"308C101C885C100C884C100C883C374C100C882C362C169C880D881C887E20CC";
		constant syscontrol_inst_instruction_ram_INIT_0A : bit_vector(0 to 255) := X"12EC882C364C173C102E191D809C10FC808C3FFC1F0C0BF0880D881C887E20CC";
		constant syscontrol_inst_instruction_ram_INIT_0B : bit_vector(0 to 255) := X"80B00BF0880D881C887E20CC300C101C885C374C100C884C362C169C883C370C";
		constant syscontrol_inst_instruction_ram_INIT_0C : bit_vector(0 to 255) := X"880C192C20CC101C887C102C100510040C701FF7880C190C887C102C0C101037";
		constant syscontrol_inst_instruction_ram_INIT_0D : bit_vector(0 to 255) := X"101C887C102C90D580C4108CCE90B05EA04F102F103E88348825100D0D101FF7";
		constant syscontrol_inst_instruction_ram_INIT_0E : bit_vector(0 to 255) := X"A0C8101C4F20A08C100C0EA010670E801FF7880C193C885C108C884C100C20CC";
		constant syscontrol_inst_instruction_ram_INIT_0F : bit_vector(0 to 255) := X"0FF050B0A00C100C0FB01077880C194C20CC101C887C102C0F3010470F101057";
		constant syscontrol_inst_instruction_ram_INIT_10 : bit_vector(0 to 255) := X"1087880C131C887C104C10A010901080100710105090A00C101C5060A00C100C";
		constant syscontrol_inst_instruction_ram_INIT_11 : bit_vector(0 to 255) := X"4D20A07C104C4C80A07C103C4750A07C101C4C20A07C100C4FC0A07C107C1100";
		constant syscontrol_inst_instruction_ram_INIT_12 : bit_vector(0 to 255) := X"808C0B3C809C0A2C12B080BC12905000A07C108C4F40A07C106C4EB0A07C105C";
		constant syscontrol_inst_instruction_ram_INIT_13 : bit_vector(0 to 255) := X"10170B3113D0880E120E887E091E884C032C883C002C882C000C881D001D1300";
		constant syscontrol_inst_instruction_ram_INIT_14 : bit_vector(0 to 255) := X"0C420B3314D0880C122C884C053C883C052C882C051C881C050C887C091C1400";
		constant syscontrol_inst_instruction_ram_INIT_15 : bit_vector(0 to 255) := X"0B3C15E0880E121E887E091E884E10BE801B883D40CD840C881C0A2C15101047";
		constant syscontrol_inst_instruction_ram_INIT_16 : bit_vector(0 to 255) := X"882C881C100C887C091C16A01057106880C080AC0E6C80AC0D5C80AC0C4C80AC";
		constant syscontrol_inst_instruction_ram_INIT_17 : bit_vector(0 to 255) := X"0B3C80AC0A2C80DC17B0880A887C091C80CC1760880C109C885C0E6C884C883C";
		constant syscontrol_inst_instruction_ram_INIT_18 : bit_vector(0 to 255) := X"000000000000000000000000000018808809887C091C80AC0D5C80AC0C4C80AC";
		constant syscontrol_inst_instruction_ram_INIT_19 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_1F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_20 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_21 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_22 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_23 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_24 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_25 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_26 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_27 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_28 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_29 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_2F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_30 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_31 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_32 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_33 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_34 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_35 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_36 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_37 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_38 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_39 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3A : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3B : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3C : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3D : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3E : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INIT_3F : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_00 : bit_vector(0 to 255) := X"EE5249EAEEEEEEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBAEBA";
		constant syscontrol_inst_instruction_ram_INITP_01 : bit_vector(0 to 255) := X"526E0E662499BBB8382403E6E0EA6EE6DFC8EBAEBAAEE9FC8EEEBAFC8EBAEBAA";
		constant syscontrol_inst_instruction_ram_INITP_02 : bit_vector(0 to 255) := X"337CDECFFB1AF3331ECCBEC607BFFFF187B3FFFDCC75249249249249BB95A492";
		constant syscontrol_inst_instruction_ram_INITP_03 : bit_vector(0 to 255) := X"000000000000000000000000000000000000000000000000000000000001F333";
		constant syscontrol_inst_instruction_ram_INITP_04 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_05 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_06 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
		constant syscontrol_inst_instruction_ram_INITP_07 : bit_vector(0 to 255) := X"0000000000000000000000000000000000000000000000000000000000000000";
